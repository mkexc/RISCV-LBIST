library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity tb_SPACE_COMP is
end entity tb_SPACE_COMP;

architecture rtl of tb_SPACE_COMP is
    component SPACE_COMP is
        port (
            D_in : in std_logic_vector(230 downto 0);
            D_out: out std_logic_vector(63 downto 0)
        );
    end component SPACE_COMP;

    signal D_in_s: std_logic_vector(230 downto 0);
    signal D_out_s: std_logic_vector(63 downto 0);

begin

    dut: SPACE_COMP
    port map (
        D_in=>D_in_s,
        D_out=>D_out_s
    );
    
   test_vect: process
   begin
        D_in_s<="100100101010101001011010010101001010101001010101001011011001010101010101010101010100010101010101100101010101010010101010101100100101010101001010101001010101010010101001010101001010101001011010010101010101100101010101010010101010101";
        wait for 10 ns;
        D_in_s<="100100101010101001011010010101001010101001010101001011011001010101010101010101010100010010101001010100101001010010101010101100100101010101001010101001010101010010101001010101001010101001011010010101010101100101010101010010101010101";
        wait for 10 ns;
        D_in_s<="100100101010101001011010010101001010101001010101001011011010010010101001010100101010010101001010000010010101000000100101010010101001010101010000100101010101111111101010100001001010101001011010010101010101100101010101010010101010101";
        wait for 10 ns;
        
        wait;
   end process test_vect;
    
    
end architecture rtl;