package CONSTANTS is
    constant N_MISR: integer := 64;
    constant N_LFSR: integer := 64;
end package CONSTANTS;