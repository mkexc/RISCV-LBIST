package constants;

parameter n_misr = 64;
parameter n_lfsr = 64;

endpackage