library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.constants.all;

entity ROM is
    port (
        addr: in std_logic_vector(3 downto 0);
        dout: out std_logic_vector(N_LFSR-1 downto 0)
    );
end entity ROM;

architecture rtl of ROM is
    type ROM_Type is array(15 downto 0) of std_logic_vector(N_LFSR-1 downto 0);
    signal rom : ROM_Type := (  0 => "1010101010101010101010101010101010101010101010101010101010101001",
                                1 => "0100100101010000100101010100101010100001001010010101001000010001",
                                2 => "1110100101010010111111110100101010101011110100000000000101010010",
                                3 => "1111111111111000000000000000111011100100111111110100100101010010",
                                4 => "0010010101001010100101111110101010100101010010000000101010101010",
                                5 => "0101010010000000000001010101111111010010101010101010100101010101",
                                6 => "1001010100000010101010100000101010010101010101010101010001010100",
                                7 => "0010101111110100101010101010010001001010101010101000101010101010",
                                8 => "1111101010101100101010101010101010100101010101000000000000011101",
                                9 => "0000000000001001010101111111010000000000010100100101000000110101",
                                10=> "0010101010101010100010010000101111101001010000010100010000010010",
                                11=> "0101010101010101001000111111111111111111111111110000000000111111",
                                others=>(N_LFSR-1 downto 0 => '0')
                                );
begin
    
    dout<=rom(to_integer(unsigned(addr)));
    
end architecture rtl;